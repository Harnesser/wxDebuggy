module feedback_1
  (
    input in1,
    output out1
  );

  two_in_two_out U1 ( .in1(in1), .in2(n2), .out1(out1), .out2(n2) );

endmodule

