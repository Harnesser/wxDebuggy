module one_in_one_out
  (
   input in,
   output out
   );
   
   
endmodule
   
