module a
  (
   input in1,
   input in2,
   output out1,
   output out2
   );
   
   
endmodule
   