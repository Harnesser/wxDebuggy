module one_in_two_out
  (
   input in,
   output out1,
   output out2
   );
   
   
endmodule
   
