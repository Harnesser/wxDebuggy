module three_in_three_out
  (
   input in1,
   input in2,
   input in3,
   output out1,
   output out2,
   output out3
   );
   
   
endmodule
   
