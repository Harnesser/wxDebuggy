module b
 ( input in1, 
   input in2,
   input in3,
   output out1,
   output out2 );
   
endmodule
   