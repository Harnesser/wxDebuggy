module two_in_three_out
  (
   input in1,
   input in2,
   output out1,
   output out2,
   output out3
   );
   
   
endmodule
   
