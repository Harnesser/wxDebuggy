module a_clk_rstb
  (
   input in1,
   input in2,
   input clk,
   input rstb,
   output out1,
   output out2
   );
   
   
endmodule
   
