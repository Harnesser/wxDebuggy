module four_in_four_out
  (
   input in1,
   input in2,
   input in3,
   input in4,
   output out1,
   output out2,
   output out3,
   output out4
   );
   
   
endmodule
   
