//
// A Simple Module declaration
//
// $Id: all_one_line.v,v 1.1 2007-08-15 23:47:37 marty Exp $

module all_one_line(input resetb,input mclk,input [3:0] din,output [6:0] dout,output do_something); endmodule // ports_only
