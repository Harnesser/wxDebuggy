module three_in_one_out
  (
   input in1,
   input in2,
   input in3,
   output out
   );
   
   
endmodule
   
