module b_clk_rstb
 ( input in1, 
   input in2,
   input in3,
   input clk,
   input rstb,
   output out1,
   output out2,
   output out3 );
   
endmodule
   
