module one_in_three_out
  (
   input in,
   output out1,
   output out2,
   output out3
   );
   
endmodule
   
