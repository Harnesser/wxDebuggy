module and2
  (
   input A,
   input B,
   output Y
   );
   
   
endmodule
   
