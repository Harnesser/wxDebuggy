module two_in
  (
   input in1,
   input in2
   );
   
   
endmodule
