module inv
  (
   input A,
   output Y
   );
   
   
endmodule
   
