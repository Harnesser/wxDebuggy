module one_in_four_out
  (
   input in1,
   output out1,
   output out2,
   output out3,
   output out4
   );
   
   
endmodule
   
