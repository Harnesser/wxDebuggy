module four_out
  (
   output out1,
   output out2,
   output out3,
   output out4
   );
   
   
endmodule
   
