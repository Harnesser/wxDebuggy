module two_in_two_out
  (
   input in1,
   input in2,
   output out1,
   output out2
   );
   
   
endmodule
   
