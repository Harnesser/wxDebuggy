module two_in_one_out
  (
   input in1,
   input in2,
   output out
   );
   
   
endmodule
   
